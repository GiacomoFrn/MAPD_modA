-- Buttons

-- Switches

-- RGB LEDs